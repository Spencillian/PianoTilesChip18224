`default_nettype none

module 
